*SAR Logic

V1 COMP 0 PULSE(0 1.8 1ns 1ns 1ns 1us 2us)
V2 RESET 0 PULSE(0 1.8 1ns 1ns 1ns .05us 6us)
V3 CLK 0 PULSE(0 1.8 1ns 1ns 1ns .25us .5us)
V5 VDD 0 1.8
X1 VDD 0 RESET CLK COMP D9 D8 D7 D6 D5 D4 D3 D2 D1 D0 EOC SAR

.include SAR.lib
.include osu018.lib
.tran 1ns 15us

.control
run
plot  V(CLK)  V(RESET)+2  V(COMP)+4
plot  V(EOC)  V(D9)+2  V(D8)+4  V(D7)+6  V(D6)+8  V(D5)+10   V(D4)+12  V(D3)+14  V(D2)+16  V(D1)+18   V(D0)+20 
.endc
.end
